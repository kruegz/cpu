package my_testbench_pkg;
  import uvm_pkg::*;
  
  `include "my_sequence.svh"
  `include "my_driver.svh"
  `include "my_agent.sv"
  `include "my_env.sv"
  `include "my_test.sv"
  
endpackage